`timescale 1ns / 1ps
/*--  *******************************************************
--  Computer Architecture Course, Laboratory Sources 
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce[dot]aut[dot]ac[dot]ir
--  *******************************************************
--  All Rights reserved (C) 2021-2022
--  *******************
--  Student ID  : 9931103
--  Student Name: Sarvin Nami
--  Student Mail: srvn0nm@gmail.com
--  *******************
--  *******************
--  Student ID  : 9931071
--  Student Name: Abtin Zandi
--  Student Mail: abtin81@aut.ac.ir
--  *******************
--  Additional Comments:
--
--*/

/*-----------------------------------------------------------
---  Module Name: adderSubtractor
-----------------------------------------------------------*/
module adderSubtractor(time_out,time_in, cin, cout, sum);
input time_out;
input time_in;
input cin;
output cout;
output sum;
 
 	 wire newTime_in;
	 xor (newTime_in, 1'b1, time_in);
	 fullAdder f(time_out,newTime_in, cin, cout, sum);

endmodule
